//`define DSP_FULL_ON
`define DSP_FULL_ON
`define USE_DSP (* USE_DSP48 = "YES" *)